module instatiate((KEY,LEDR,SW,HEX0,HEX1,HEX2,HEX3);